module shift(
  clock,
  data_in,
  data_out
);
	parameter width=10;
	
	input clock;
	input      [width-1:0] data_in;
	output reg [width-1:0] data_out;
 
	always @(posedge clock) data_out <= data_in;
	
 endmodule