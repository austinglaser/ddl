module fir(
  clock,
  data_in,
  data_out
);
  //parameters
	parameter width =  10;
	parameter length = 465;
	parameter n_coeffs = 465;
	parameter ones = 0;
	
	// define arguments
	input clock;
	input  [width-1:0] data_in;
	output [width-1:0] data_out;
	
	// two-dimensional coefficient registers (initialized in 'initial' block)
	reg [16:0] coeff [n_coeffs-1:0];
	
	// 
	wire [width-1:0] 			data_values [length-1:0];
	wire [(width + 17)-1:0]	mult_values [length-1:0];
	wire [(width + 17)-1:0]	sum_values  [length-1:0];
	
	assign data_out = sum_values[length-1] >> 15;
	
	shift_reg #(width, length) data_shift(clock, data_in, data_values);
	
	assign sum_values[0]  = mult_values[0];
	
	genvar i;
	generate
		for (i = 0; i < length; i = i+1) begin:fir_gen
			multiply #(width, 17) MULT(clock, data_values[i], coeff[(n_coeffs-1)-i], mult_values[i]);
			
			if (i == 0) assign sum_values[i] = mult_values[i];
			else			assign sum_values[i] = mult_values[i] + sum_values[i-1];
		end
	endgenerate
	
	initial begin
  		coeff[0]   =  17'd442;	// This coefficient should be multiplied with the oldest input value
  		coeff[1]   = -17'd373;
  		coeff[2]   = -17'd169;
  		coeff[3]   = -17'd37;
  		coeff[4]   =  17'd20;
  		coeff[5]   =  17'd15;
  		coeff[6]   = -17'd21;
  		coeff[7]   = -17'd61;
  		coeff[8]   = -17'd80;
  		coeff[9]   = -17'd70;
  		coeff[10]  = -17'd37;
  		coeff[11]  =  17'd4;
  		coeff[12]  =  17'd35;
  		coeff[13]  =  17'd45;
  		coeff[14]  =  17'd32;
  		coeff[15]  =  17'd3;
  		coeff[16]  = -17'd29;
  		coeff[17]  = -17'd49;
  		coeff[18]  = -17'd49;
  		coeff[19]  = -17'd30;
  		coeff[20]  =  17'd0;
  		coeff[21]  =  17'd29;
  		coeff[22]  =  17'd44;
  		coeff[23]  =  17'd41;
  		coeff[24]  =  17'd22;
  		coeff[25]  = -17'd6;
  		coeff[26]  = -17'd31;
  		coeff[27]  = -17'd43;
  		coeff[28]  = -17'd37;
  		coeff[29]  = -17'd18;
  		coeff[30]  =  17'd8;
  		coeff[31]  =  17'd29;
  		coeff[32]  =  17'd38;
  		coeff[33]  =  17'd31;
  		coeff[34]  =  17'd13;
  		coeff[35]  = -17'd9;
  		coeff[36]  = -17'd25;
  		coeff[37]  = -17'd31;
  		coeff[38]  = -17'd24;
  		coeff[39]  = -17'd9;
  		coeff[40]  =  17'd8;
  		coeff[41]  =  17'd19;
  		coeff[42]  =  17'd21;
  		coeff[43]  =  17'd15;
  		coeff[44]  =  17'd4;
  		coeff[45]  = -17'd6;
  		coeff[46]  = -17'd11;
  		coeff[47]  = -17'd10;
  		coeff[48]  = -17'd4;
  		coeff[49]  =  17'd1;
  		coeff[50]  =  17'd3;
  		coeff[51]  =  17'd1;
  		coeff[52]  = -17'd4;
  		coeff[53]  = -17'd7;
  		coeff[54]  = -17'd7;
  		coeff[55]  = -17'd1;
  		coeff[56]  =  17'd10;
  		coeff[57]  =  17'd19;
  		coeff[58]  =  17'd21;
  		coeff[59]  =  17'd13;
  		coeff[60]  = -17'd3;
  		coeff[61]  = -17'd21;
  		coeff[62]  = -17'd34;
  		coeff[63]  = -17'd34;
  		coeff[64]  = -17'd19;
  		coeff[65]  =  17'd7;
  		coeff[66]  =  17'd33;
  		coeff[67]  =  17'd49;
  		coeff[68]  =  17'd47;
  		coeff[69]  =  17'd25;
  		coeff[70]  = -17'd10;
  		coeff[71]  = -17'd44;
  		coeff[72]  = -17'd63;
  		coeff[73]  = -17'd58;
  		coeff[74]  = -17'd29;
  		coeff[75]  =  17'd13;
  		coeff[76]  =  17'd52;
  		coeff[77]  =  17'd73;
  		coeff[78]  =  17'd66;
  		coeff[79]  =  17'd33;
  		coeff[80]  = -17'd15;
  		coeff[81]  = -17'd58;
  		coeff[82]  = -17'd80;
  		coeff[83]  = -17'd70;
  		coeff[84]  = -17'd34;
  		coeff[85]  =  17'd16;
  		coeff[86]  =  17'd60;
  		coeff[87]  =  17'd80;
  		coeff[88]  =  17'd69;
  		coeff[89]  =  17'd32;
  		coeff[90]  = -17'd16;
  		coeff[91]  = -17'd57;
  		coeff[92]  = -17'd75;
  		coeff[93]  = -17'd63;
  		coeff[94]  = -17'd29;
  		coeff[95]  =  17'd15;
  		coeff[96]  =  17'd50;
  		coeff[97]  =  17'd63;
  		coeff[98]  =  17'd51;
  		coeff[99]  =  17'd22;
  		coeff[100] = -17'd12;
  		coeff[101] = -17'd37;
  		coeff[102] = -17'd44;
  		coeff[103] = -17'd34;
  		coeff[104] = -17'd13;
  		coeff[105] =  17'd7;
  		coeff[106] =  17'd19;
  		coeff[107] =  17'd19;
  		coeff[108] =  17'd11;
  		coeff[109] =  17'd2;
  		coeff[110] = -17'd1;
  		coeff[111] =  17'd3;
  		coeff[112] =  17'd11;
  		coeff[113] =  17'd16;
  		coeff[114] =  17'd10;
  		coeff[115] = -17'd7;
  		coeff[116] = -17'd29;
  		coeff[117] = -17'd46;
  		coeff[118] = -17'd46;
  		coeff[119] = -17'd24;
  		coeff[120] =  17'd15;
  		coeff[121] =  17'd56;
  		coeff[122] =  17'd81;
  		coeff[123] =  17'd76;
  		coeff[124] =  17'd37;
  		coeff[125] = -17'd24;
  		coeff[126] = -17'd83;
  		coeff[127] = -17'd116;
  		coeff[128] = -17'd105;
  		coeff[129] = -17'd50;
  		coeff[130] =  17'd32;
  		coeff[131] =  17'd109;
  		coeff[132] =  17'd148;
  		coeff[133] =  17'd131;
  		coeff[134] =  17'd60;
  		coeff[135] = -17'd39;
  		coeff[136] = -17'd130;
  		coeff[137] = -17'd173;
  		coeff[138] = -17'd151;
  		coeff[139] = -17'd68;
  		coeff[140] =  17'd45;
  		coeff[141] =  17'd144;
  		coeff[142] =  17'd190;
  		coeff[143] =  17'd162;
  		coeff[144] =  17'd71;
  		coeff[145] = -17'd48;
  		coeff[146] = -17'd150;
  		coeff[147] = -17'd194;
  		coeff[148] = -17'd163;
  		coeff[149] = -17'd70;
  		coeff[150] =  17'd48;
  		coeff[151] =  17'd145;
  		coeff[152] =  17'd184;
  		coeff[153] =  17'd152;
  		coeff[154] =  17'd64;
  		coeff[155] = -17'd44;
  		coeff[156] = -17'd128;
  		coeff[157] = -17'd159;
  		coeff[158] = -17'd127;
  		coeff[159] = -17'd51;
  		coeff[160] =  17'd35;
  		coeff[161] =  17'd98;
  		coeff[162] =  17'd116;
  		coeff[163] =  17'd88;
  		coeff[164] =  17'd33;
  		coeff[165] = -17'd22;
  		coeff[166] = -17'd55;
  		coeff[167] = -17'd57;
  		coeff[168] = -17'd36;
  		coeff[169] = -17'd10;
  		coeff[170] =  17'd4;
  		coeff[171] = -17'd2;
  		coeff[172] = -17'd19;
  		coeff[173] = -17'd30;
  		coeff[174] = -17'd19;
  		coeff[175] =  17'd19;
  		coeff[176] =  17'd71;
  		coeff[177] =  17'd110;
  		coeff[178] =  17'd108;
  		coeff[179] =  17'd52;
  		coeff[180] = -17'd47;
  		coeff[181] = -17'd151;
  		coeff[182] = -17'd214;
  		coeff[183] = -17'd196;
  		coeff[184] = -17'd88;
  		coeff[185] =  17'd78;
  		coeff[186] =  17'd240;
  		coeff[187] =  17'd327;
  		coeff[188] =  17'd290;
  		coeff[189] =  17'd126;
  		coeff[190] = -17'd111;
  		coeff[191] = -17'd333;
  		coeff[192] = -17'd445;
  		coeff[193] = -17'd387;
  		coeff[194] = -17'd165;
  		coeff[195] =  17'd147;
  		coeff[196] =  17'd429;
  		coeff[197] =  17'd564;
  		coeff[198] =  17'd484;
  		coeff[199] =  17'd202;
  		coeff[200] = -17'd183;
  		coeff[201] = -17'd523;
  		coeff[202] = -17'd680;
  		coeff[203] = -17'd577;
  		coeff[204] = -17'd237;
  		coeff[205] =  17'd217;
  		coeff[206] =  17'd613;
  		coeff[207] =  17'd788;
  		coeff[208] =  17'd662;
  		coeff[209] =  17'd269;
  		coeff[210] = -17'd249;
  		coeff[211] = -17'd693;
  		coeff[212] = -17'd883;
  		coeff[213] = -17'd736;
  		coeff[214] = -17'd294;
  		coeff[215] =  17'd278;
  		coeff[216] =  17'd761;
  		coeff[217] =  17'd962;
  		coeff[218] =  17'd795;
  		coeff[219] =  17'd314;
  		coeff[220] = -17'd301;
  		coeff[221] = -17'd813;
  		coeff[222] = -17'd1021;
  		coeff[223] = -17'd837;
  		coeff[224] = -17'd326;
  		coeff[225] =  17'd318;
  		coeff[226] =  17'd848;
  		coeff[227] =  17'd1057;
  		coeff[228] =  17'd861;
  		coeff[229] =  17'd331;
  		coeff[230] = -17'd329;
  		coeff[231] = -17'd865;
  		coeff[232] =  17'd31698;
  		coeff[233] = -17'd865;
  		coeff[234] = -17'd329;
  		coeff[235] =  17'd331;
  		coeff[236] =  17'd861;
  		coeff[237] =  17'd1057;
  		coeff[238] =  17'd848;
  		coeff[239] =  17'd318;
  		coeff[240] = -17'd326;
  		coeff[241] = -17'd837;
  		coeff[242] = -17'd1021;
  		coeff[243] = -17'd813;
  		coeff[244] = -17'd301;
  		coeff[245] =  17'd314;
  		coeff[246] =  17'd795;
  		coeff[247] =  17'd962;
  		coeff[248] =  17'd761;
  		coeff[249] =  17'd278;
  		coeff[250] = -17'd294;
  		coeff[251] = -17'd736;
  		coeff[252] = -17'd883;
  		coeff[253] = -17'd693;
  		coeff[254] = -17'd249;
  		coeff[255] =  17'd269;
  		coeff[256] =  17'd662;
  		coeff[257] =  17'd788;
  		coeff[258] =  17'd613;
  		coeff[259] =  17'd217;
  		coeff[260] = -17'd237;
  		coeff[261] = -17'd577;
  		coeff[262] = -17'd680;
  		coeff[263] = -17'd523;
  		coeff[264] = -17'd183;
  		coeff[265] =  17'd202;
  		coeff[266] =  17'd484;
  		coeff[267] =  17'd564;
  		coeff[268] =  17'd429;
  		coeff[269] =  17'd147;
  		coeff[270] = -17'd165;
  		coeff[271] = -17'd387;
  		coeff[272] = -17'd445;
  		coeff[273] = -17'd333;
  		coeff[274] = -17'd111;
  		coeff[275] =  17'd126;
  		coeff[276] =  17'd290;
  		coeff[277] =  17'd327;
  		coeff[278] =  17'd240;
  		coeff[279] =  17'd78;
  		coeff[280] = -17'd88;
  		coeff[281] = -17'd196;
  		coeff[282] = -17'd214;
  		coeff[283] = -17'd151;
  		coeff[284] = -17'd47;
  		coeff[285] =  17'd52;
  		coeff[286] =  17'd108;
  		coeff[287] =  17'd110;
  		coeff[288] =  17'd71;
  		coeff[289] =  17'd19;
  		coeff[290] = -17'd19;
  		coeff[291] = -17'd30;
  		coeff[292] = -17'd19;
  		coeff[293] = -17'd2;
  		coeff[294] =  17'd4;
  		coeff[295] = -17'd10;
  		coeff[296] = -17'd36;
  		coeff[297] = -17'd57;
  		coeff[298] = -17'd55;
  		coeff[299] = -17'd22;
  		coeff[300] =  17'd33;
  		coeff[301] =  17'd88;
  		coeff[302] =  17'd116;
  		coeff[303] =  17'd98;
  		coeff[304] =  17'd35;
  		coeff[305] = -17'd51;
  		coeff[306] = -17'd127;
  		coeff[307] = -17'd159;
  		coeff[308] = -17'd128;
  		coeff[309] = -17'd44;
  		coeff[310] =  17'd64;
  		coeff[311] =  17'd152;
  		coeff[312] =  17'd184;
  		coeff[313] =  17'd145;
  		coeff[314] =  17'd48;
  		coeff[315] = -17'd70;
  		coeff[316] = -17'd163;
  		coeff[317] = -17'd194;
  		coeff[318] = -17'd150;
  		coeff[319] = -17'd48;
  		coeff[320] =  17'd71;
  		coeff[321] =  17'd162;
  		coeff[322] =  17'd190;
  		coeff[323] =  17'd144;
  		coeff[324] =  17'd45;
  		coeff[325] = -17'd68;
  		coeff[326] = -17'd151;
  		coeff[327] = -17'd173;
  		coeff[328] = -17'd130;
  		coeff[329] = -17'd39;
  		coeff[330] =  17'd60;
  		coeff[331] =  17'd131;
  		coeff[332] =  17'd148;
  		coeff[333] =  17'd109;
  		coeff[334] =  17'd32;
  		coeff[335] = -17'd50;
  		coeff[336] = -17'd105;
  		coeff[337] = -17'd116;
  		coeff[338] = -17'd83;
  		coeff[339] = -17'd24;
  		coeff[340] =  17'd37;
  		coeff[341] =  17'd76;
  		coeff[342] =  17'd81;
  		coeff[343] =  17'd56;
  		coeff[344] =  17'd15;
  		coeff[345] = -17'd24;
  		coeff[346] = -17'd46;
  		coeff[347] = -17'd46;
  		coeff[348] = -17'd29;
  		coeff[349] = -17'd7;
  		coeff[350] =  17'd10;
  		coeff[351] =  17'd16;
  		coeff[352] =  17'd11;
  		coeff[353] =  17'd3;
  		coeff[354] = -17'd1;
  		coeff[355] =  17'd2;
  		coeff[356] =  17'd11;
  		coeff[357] =  17'd19;
  		coeff[358] =  17'd19;
  		coeff[359] =  17'd7;
  		coeff[360] = -17'd13;
  		coeff[361] = -17'd34;
  		coeff[362] = -17'd44;
  		coeff[363] = -17'd37;
  		coeff[364] = -17'd12;
  		coeff[365] =  17'd22;
  		coeff[366] =  17'd51;
  		coeff[367] =  17'd63;
  		coeff[368] =  17'd50;
  		coeff[369] =  17'd15;
  		coeff[370] = -17'd29;
  		coeff[371] = -17'd63;
  		coeff[372] = -17'd75;
  		coeff[373] = -17'd57;
  		coeff[374] = -17'd16;
  		coeff[375] =  17'd32;
  		coeff[376] =  17'd69;
  		coeff[377] =  17'd80;
  		coeff[378] =  17'd60;
  		coeff[379] =  17'd16;
  		coeff[380] = -17'd34;
  		coeff[381] = -17'd70;
  		coeff[382] = -17'd80;
  		coeff[383] = -17'd58;
  		coeff[384] = -17'd15;
  		coeff[385] =  17'd33;
  		coeff[386] =  17'd66;
  		coeff[387] =  17'd73;
  		coeff[388] =  17'd52;
  		coeff[389] =  17'd13;
  		coeff[390] = -17'd29;
  		coeff[391] = -17'd58;
  		coeff[392] = -17'd63;
  		coeff[393] = -17'd44;
  		coeff[394] = -17'd10;
  		coeff[395] =  17'd25;
  		coeff[396] =  17'd47;
  		coeff[397] =  17'd49;
  		coeff[398] =  17'd33;
  		coeff[399] =  17'd7;
  		coeff[400] = -17'd19;
  		coeff[401] = -17'd34;
  		coeff[402] = -17'd34;
  		coeff[403] = -17'd21;
  		coeff[404] = -17'd3;
  		coeff[405] =  17'd13;
  		coeff[406] =  17'd21;
  		coeff[407] =  17'd19;
  		coeff[408] =  17'd10;
  		coeff[409] = -17'd1;
  		coeff[410] = -17'd7;
  		coeff[411] = -17'd7;
  		coeff[412] = -17'd4;
  		coeff[413] =  17'd1;
  		coeff[414] =  17'd3;
  		coeff[415] =  17'd1;
  		coeff[416] = -17'd4;
  		coeff[417] = -17'd10;
  		coeff[418] = -17'd11;
  		coeff[419] = -17'd6;
  		coeff[420] =  17'd4;
  		coeff[421] =  17'd15;
  		coeff[422] =  17'd21;
  		coeff[423] =  17'd19;
  		coeff[424] =  17'd8;
  		coeff[425] = -17'd9;
  		coeff[426] = -17'd24;
  		coeff[427] = -17'd31;
  		coeff[428] = -17'd25;
  		coeff[429] = -17'd9;
  		coeff[430] =  17'd13;
  		coeff[431] =  17'd31;
  		coeff[432] =  17'd38;
  		coeff[433] =  17'd29;
  		coeff[434] =  17'd8;
  		coeff[435] = -17'd18;
  		coeff[436] = -17'd37;
  		coeff[437] = -17'd43;
  		coeff[438] = -17'd31;
  		coeff[439] = -17'd6;
  		coeff[440] =  17'd22;
  		coeff[441] =  17'd41;
  		coeff[442] =  17'd44;
  		coeff[443] =  17'd29;
  		coeff[444] =  17'd0;
  		coeff[445] = -17'd30;
  		coeff[446] = -17'd49;
  		coeff[447] = -17'd49;
  		coeff[448] = -17'd29;
  		coeff[449] =  17'd3;
  		coeff[450] =  17'd32;
  		coeff[451] =  17'd45;
  		coeff[452] =  17'd35;
  		coeff[453] =  17'd4;
  		coeff[454] = -17'd37;
  		coeff[455] = -17'd70;
  		coeff[456] = -17'd80;
  		coeff[457] = -17'd61;
  		coeff[458] = -17'd21;
  		coeff[459] =  17'd15;
  		coeff[460] =  17'd20;
  		coeff[461] = -17'd37;
  		coeff[462] = -17'd169;
  		coeff[463] = -17'd373;
  		coeff[464] =  17'd442;
	end

endmodule
