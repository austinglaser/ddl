library verilog;
use verilog.vl_types.all;
entity mux6 is
    generic(
        width           : integer := 1
    );
    port(
        d0              : in     vl_logic_vector;
        d1              : in     vl_logic_vector;
        d2              : in     vl_logic_vector;
        d3              : in     vl_logic_vector;
        d4              : in     vl_logic_vector;
        d5              : in     vl_logic_vector;
        s               : in     vl_logic_vector(2 downto 0);
        y               : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of width : constant is 1;
end mux6;
