module coeff_calc (
    coeff
);
  // parameters define which coefficient this will have
  parameter coeffIndex = 0;
  parameter ones = 0;
  
  // define argument
  output reg [16:0] coeff;
  
  always @ (*) begin
    if (ones) coeff = 17'd1; // for debug purposes
    else
      case ( coeffIndex )
      
        12'd0: coeff   =  17'd442; // This coefficient should be multiplied with the oldest input value
        12'd1: coeff   = -17'd373;
        12'd2: coeff   = -17'd169;
        12'd3: coeff   = -17'd37;
        12'd4: coeff   =  17'd20;
        12'd5: coeff   =  17'd15;
        12'd6: coeff   = -17'd21;
        12'd7: coeff   = -17'd61;
        12'd8: coeff   = -17'd80;
        12'd9: coeff   = -17'd70;
        12'd10: coeff  = -17'd37;
        12'd11: coeff  =  17'd4;
        12'd12: coeff  =  17'd35;
        12'd13: coeff  =  17'd45;
        12'd14: coeff  =  17'd32;
        12'd15: coeff  =  17'd3;
        12'd16: coeff  = -17'd29;
        12'd17: coeff  = -17'd49;
        12'd18: coeff  = -17'd49;
        12'd19: coeff  = -17'd30;
        12'd20: coeff  =  17'd0;
        12'd21: coeff  =  17'd29;
        12'd22: coeff  =  17'd44;
        12'd23: coeff  =  17'd41;
        12'd24: coeff  =  17'd22;
        12'd25: coeff  = -17'd6;
        12'd26: coeff  = -17'd31;
        12'd27: coeff  = -17'd43;
        12'd28: coeff  = -17'd37;
        12'd29: coeff  = -17'd18;
        12'd30: coeff  =  17'd8;
        12'd31: coeff  =  17'd29;
        12'd32: coeff  =  17'd38;
        12'd33: coeff  =  17'd31;
        12'd34: coeff  =  17'd13;
        12'd35: coeff  = -17'd9;
        12'd36: coeff  = -17'd25;
        12'd37: coeff  = -17'd31;
        12'd38: coeff  = -17'd24;
        12'd39: coeff  = -17'd9;
        12'd40: coeff  =  17'd8;
        12'd41: coeff  =  17'd19;
        12'd42: coeff  =  17'd21;
        12'd43: coeff  =  17'd15;
        12'd44: coeff  =  17'd4;
        12'd45: coeff  = -17'd6;
        12'd46: coeff  = -17'd11;
        12'd47: coeff  = -17'd10;
        12'd48: coeff  = -17'd4;
        12'd49: coeff  =  17'd1;
        12'd50: coeff  =  17'd3;
        12'd51: coeff  =  17'd1;
        12'd52: coeff  = -17'd4;
        12'd53: coeff  = -17'd7;
        12'd54: coeff  = -17'd7;
        12'd55: coeff  = -17'd1;
        12'd56: coeff  =  17'd10;
        12'd57: coeff  =  17'd19;
        12'd58: coeff  =  17'd21;
        12'd59: coeff  =  17'd13;
        12'd60: coeff  = -17'd3;
        12'd61: coeff  = -17'd21;
        12'd62: coeff  = -17'd34;
        12'd63: coeff  = -17'd34;
        12'd64: coeff  = -17'd19;
        12'd65: coeff  =  17'd7;
        12'd66: coeff  =  17'd33;
        12'd67: coeff  =  17'd49;
        12'd68: coeff  =  17'd47;
        12'd69: coeff  =  17'd25;
        12'd70: coeff  = -17'd10;
        12'd71: coeff  = -17'd44;
        12'd72: coeff  = -17'd63;
        12'd73: coeff  = -17'd58;
        12'd74: coeff  = -17'd29;
        12'd75: coeff  =  17'd13;
        12'd76: coeff  =  17'd52;
        12'd77: coeff  =  17'd73;
        12'd78: coeff  =  17'd66;
        12'd79: coeff  =  17'd33;
        12'd80: coeff  = -17'd15;
        12'd81: coeff  = -17'd58;
        12'd82: coeff  = -17'd80;
        12'd83: coeff  = -17'd70;
        12'd84: coeff  = -17'd34;
        12'd85: coeff  =  17'd16;
        12'd86: coeff  =  17'd60;
        12'd87: coeff  =  17'd80;
        12'd88: coeff  =  17'd69;
        12'd89: coeff  =  17'd32;
        12'd90: coeff  = -17'd16;
        12'd91: coeff  = -17'd57;
        12'd92: coeff  = -17'd75;
        12'd93: coeff  = -17'd63;
        12'd94: coeff  = -17'd29;
        12'd95: coeff  =  17'd15;
        12'd96: coeff  =  17'd50;
        12'd97: coeff  =  17'd63;
        12'd98: coeff  =  17'd51;
        12'd99: coeff  =  17'd22;
        12'd100: coeff = -17'd12;
        12'd101: coeff = -17'd37;
        12'd102: coeff = -17'd44;
        12'd103: coeff = -17'd34;
        12'd104: coeff = -17'd13;
        12'd105: coeff =  17'd7;
        12'd106: coeff =  17'd19;
        12'd107: coeff =  17'd19;
        12'd108: coeff =  17'd11;
        12'd109: coeff =  17'd2;
        12'd110: coeff = -17'd1;
        12'd111: coeff =  17'd3;
        12'd112: coeff =  17'd11;
        12'd113: coeff =  17'd16;
        12'd114: coeff =  17'd10;
        12'd115: coeff = -17'd7;
        12'd116: coeff = -17'd29;
        12'd117: coeff = -17'd46;
        12'd118: coeff = -17'd46;
        12'd119: coeff = -17'd24;
        12'd120: coeff =  17'd15;
        12'd121: coeff =  17'd56;
        12'd122: coeff =  17'd81;
        12'd123: coeff =  17'd76;
        12'd124: coeff =  17'd37;
        12'd125: coeff = -17'd24;
        12'd126: coeff = -17'd83;
        12'd127: coeff = -17'd116;
        12'd128: coeff = -17'd105;
        12'd129: coeff = -17'd50;
        12'd130: coeff =  17'd32;
        12'd131: coeff =  17'd109;
        12'd132: coeff =  17'd148;
        12'd133: coeff =  17'd131;
        12'd134: coeff =  17'd60;
        12'd135: coeff = -17'd39;
        12'd136: coeff = -17'd130;
        12'd137: coeff = -17'd173;
        12'd138: coeff = -17'd151;
        12'd139: coeff = -17'd68;
        12'd140: coeff =  17'd45;
        12'd141: coeff =  17'd144;
        12'd142: coeff =  17'd190;
        12'd143: coeff =  17'd162;
        12'd144: coeff =  17'd71;
        12'd145: coeff = -17'd48;
        12'd146: coeff = -17'd150;
        12'd147: coeff = -17'd194;
        12'd148: coeff = -17'd163;
        12'd149: coeff = -17'd70;
        12'd150: coeff =  17'd48;
        12'd151: coeff =  17'd145;
        12'd152: coeff =  17'd184;
        12'd153: coeff =  17'd152;
        12'd154: coeff =  17'd64;
        12'd155: coeff = -17'd44;
        12'd156: coeff = -17'd128;
        12'd157: coeff = -17'd159;
        12'd158: coeff = -17'd127;
        12'd159: coeff = -17'd51;
        12'd160: coeff =  17'd35;
        12'd161: coeff =  17'd98;
        12'd162: coeff =  17'd116;
        12'd163: coeff =  17'd88;
        12'd164: coeff =  17'd33;
        12'd165: coeff = -17'd22;
        12'd166: coeff = -17'd55;
        12'd167: coeff = -17'd57;
        12'd168: coeff = -17'd36;
        12'd169: coeff = -17'd10;
        12'd170: coeff =  17'd4;
        12'd171: coeff = -17'd2;
        12'd172: coeff = -17'd19;
        12'd173: coeff = -17'd30;
        12'd174: coeff = -17'd19;
        12'd175: coeff =  17'd19;
        12'd176: coeff =  17'd71;
        12'd177: coeff =  17'd110;
        12'd178: coeff =  17'd108;
        12'd179: coeff =  17'd52;
        12'd180: coeff = -17'd47;
        12'd181: coeff = -17'd151;
        12'd182: coeff = -17'd214;
        12'd183: coeff = -17'd196;
        12'd184: coeff = -17'd88;
        12'd185: coeff =  17'd78;
        12'd186: coeff =  17'd240;
        12'd187: coeff =  17'd327;
        12'd188: coeff =  17'd290;
        12'd189: coeff =  17'd126;
        12'd190: coeff = -17'd111;
        12'd191: coeff = -17'd333;
        12'd192: coeff = -17'd445;
        12'd193: coeff = -17'd387;
        12'd194: coeff = -17'd165;
        12'd195: coeff =  17'd147;
        12'd196: coeff =  17'd429;
        12'd197: coeff =  17'd564;
        12'd198: coeff =  17'd484;
        12'd199: coeff =  17'd202;
        12'd200: coeff = -17'd183;
        12'd201: coeff = -17'd523;
        12'd202: coeff = -17'd680;
        12'd203: coeff = -17'd577;
        12'd204: coeff = -17'd237;
        12'd205: coeff =  17'd217;
        12'd206: coeff =  17'd613;
        12'd207: coeff =  17'd788;
        12'd208: coeff =  17'd662;
        12'd209: coeff =  17'd269;
        12'd210: coeff = -17'd249;
        12'd211: coeff = -17'd693;
        12'd212: coeff = -17'd883;
        12'd213: coeff = -17'd736;
        12'd214: coeff = -17'd294;
        12'd215: coeff =  17'd278;
        12'd216: coeff =  17'd761;
        12'd217: coeff =  17'd962;
        12'd218: coeff =  17'd795;
        12'd219: coeff =  17'd314;
        12'd220: coeff = -17'd301;
        12'd221: coeff = -17'd813;
        12'd222: coeff = -17'd1021;
        12'd223: coeff = -17'd837;
        12'd224: coeff = -17'd326;
        12'd225: coeff =  17'd318;
        12'd226: coeff =  17'd848;
        12'd227: coeff =  17'd1057;
        12'd228: coeff =  17'd861;
        12'd229: coeff =  17'd331;
        12'd230: coeff = -17'd329;
        12'd231: coeff = -17'd865;
        12'd232: coeff =  17'd31698;
        12'd233: coeff = -17'd865;
        12'd234: coeff = -17'd329;
        12'd235: coeff =  17'd331;
        12'd236: coeff =  17'd861;
        12'd237: coeff =  17'd1057;
        12'd238: coeff =  17'd848;
        12'd239: coeff =  17'd318;
        12'd240: coeff = -17'd326;
        12'd241: coeff = -17'd837;
        12'd242: coeff = -17'd1021;
        12'd243: coeff = -17'd813;
        12'd244: coeff = -17'd301;
        12'd245: coeff =  17'd314;
        12'd246: coeff =  17'd795;
        12'd247: coeff =  17'd962;
        12'd248: coeff =  17'd761;
        12'd249: coeff =  17'd278;
        12'd250: coeff = -17'd294;
        12'd251: coeff = -17'd736;
        12'd252: coeff = -17'd883;
        12'd253: coeff = -17'd693;
        12'd254: coeff = -17'd249;
        12'd255: coeff =  17'd269;
        12'd256: coeff =  17'd662;
        12'd257: coeff =  17'd788;
        12'd258: coeff =  17'd613;
        12'd259: coeff =  17'd217;
        12'd260: coeff = -17'd237;
        12'd261: coeff = -17'd577;
        12'd262: coeff = -17'd680;
        12'd263: coeff = -17'd523;
        12'd264: coeff = -17'd183;
        12'd265: coeff =  17'd202;
        12'd266: coeff =  17'd484;
        12'd267: coeff =  17'd564;
        12'd268: coeff =  17'd429;
        12'd269: coeff =  17'd147;
        12'd270: coeff = -17'd165;
        12'd271: coeff = -17'd387;
        12'd272: coeff = -17'd445;
        12'd273: coeff = -17'd333;
        12'd274: coeff = -17'd111;
        12'd275: coeff =  17'd126;
        12'd276: coeff =  17'd290;
        12'd277: coeff =  17'd327;
        12'd278: coeff =  17'd240;
        12'd279: coeff =  17'd78;
        12'd280: coeff = -17'd88;
        12'd281: coeff = -17'd196;
        12'd282: coeff = -17'd214;
        12'd283: coeff = -17'd151;
        12'd284: coeff = -17'd47;
        12'd285: coeff =  17'd52;
        12'd286: coeff =  17'd108;
        12'd287: coeff =  17'd110;
        12'd288: coeff =  17'd71;
        12'd289: coeff =  17'd19;
        12'd290: coeff = -17'd19;
        12'd291: coeff = -17'd30;
        12'd292: coeff = -17'd19;
        12'd293: coeff = -17'd2;
        12'd294: coeff =  17'd4;
        12'd295: coeff = -17'd10;
        12'd296: coeff = -17'd36;
        12'd297: coeff = -17'd57;
        12'd298: coeff = -17'd55;
        12'd299: coeff = -17'd22;
        12'd300: coeff =  17'd33;
        12'd301: coeff =  17'd88;
        12'd302: coeff =  17'd116;
        12'd303: coeff =  17'd98;
        12'd304: coeff =  17'd35;
        12'd305: coeff = -17'd51;
        12'd306: coeff = -17'd127;
        12'd307: coeff = -17'd159;
        12'd308: coeff = -17'd128;
        12'd309: coeff = -17'd44;
        12'd310: coeff =  17'd64;
        12'd311: coeff =  17'd152;
        12'd312: coeff =  17'd184;
        12'd313: coeff =  17'd145;
        12'd314: coeff =  17'd48;
        12'd315: coeff = -17'd70;
        12'd316: coeff = -17'd163;
        12'd317: coeff = -17'd194;
        12'd318: coeff = -17'd150;
        12'd319: coeff = -17'd48;
        12'd320: coeff =  17'd71;
        12'd321: coeff =  17'd162;
        12'd322: coeff =  17'd190;
        12'd323: coeff =  17'd144;
        12'd324: coeff =  17'd45;
        12'd325: coeff = -17'd68;
        12'd326: coeff = -17'd151;
        12'd327: coeff = -17'd173;
        12'd328: coeff = -17'd130;
        12'd329: coeff = -17'd39;
        12'd330: coeff =  17'd60;
        12'd331: coeff =  17'd131;
        12'd332: coeff =  17'd148;
        12'd333: coeff =  17'd109;
        12'd334: coeff =  17'd32;
        12'd335: coeff = -17'd50;
        12'd336: coeff = -17'd105;
        12'd337: coeff = -17'd116;
        12'd338: coeff = -17'd83;
        12'd339: coeff = -17'd24;
        12'd340: coeff =  17'd37;
        12'd341: coeff =  17'd76;
        12'd342: coeff =  17'd81;
        12'd343: coeff =  17'd56;
        12'd344: coeff =  17'd15;
        12'd345: coeff = -17'd24;
        12'd346: coeff = -17'd46;
        12'd347: coeff = -17'd46;
        12'd348: coeff = -17'd29;
        12'd349: coeff = -17'd7;
        12'd350: coeff =  17'd10;
        12'd351: coeff =  17'd16;
        12'd352: coeff =  17'd11;
        12'd353: coeff =  17'd3;
        12'd354: coeff = -17'd1;
        12'd355: coeff =  17'd2;
        12'd356: coeff =  17'd11;
        12'd357: coeff =  17'd19;
        12'd358: coeff =  17'd19;
        12'd359: coeff =  17'd7;
        12'd360: coeff = -17'd13;
        12'd361: coeff = -17'd34;
        12'd362: coeff = -17'd44;
        12'd363: coeff = -17'd37;
        12'd364: coeff = -17'd12;
        12'd365: coeff =  17'd22;
        12'd366: coeff =  17'd51;
        12'd367: coeff =  17'd63;
        12'd368: coeff =  17'd50;
        12'd369: coeff =  17'd15;
        12'd370: coeff = -17'd29;
        12'd371: coeff = -17'd63;
        12'd372: coeff = -17'd75;
        12'd373: coeff = -17'd57;
        12'd374: coeff = -17'd16;
        12'd375: coeff =  17'd32;
        12'd376: coeff =  17'd69;
        12'd377: coeff =  17'd80;
        12'd378: coeff =  17'd60;
        12'd379: coeff =  17'd16;
        12'd380: coeff = -17'd34;
        12'd381: coeff = -17'd70;
        12'd382: coeff = -17'd80;
        12'd383: coeff = -17'd58;
        12'd384: coeff = -17'd15;
        12'd385: coeff =  17'd33;
        12'd386: coeff =  17'd66;
        12'd387: coeff =  17'd73;
        12'd388: coeff =  17'd52;
        12'd389: coeff =  17'd13;
        12'd390: coeff = -17'd29;
        12'd391: coeff = -17'd58;
        12'd392: coeff = -17'd63;
        12'd393: coeff = -17'd44;
        12'd394: coeff = -17'd10;
        12'd395: coeff =  17'd25;
        12'd396: coeff =  17'd47;
        12'd397: coeff =  17'd49;
        12'd398: coeff =  17'd33;
        12'd399: coeff =  17'd7;
        12'd400: coeff = -17'd19;
        12'd401: coeff = -17'd34;
        12'd402: coeff = -17'd34;
        12'd403: coeff = -17'd21;
        12'd404: coeff = -17'd3;
        12'd405: coeff =  17'd13;
        12'd406: coeff =  17'd21;
        12'd407: coeff =  17'd19;
        12'd408: coeff =  17'd10;
        12'd409: coeff = -17'd1;
        12'd410: coeff = -17'd7;
        12'd411: coeff = -17'd7;
        12'd412: coeff = -17'd4;
        12'd413: coeff =  17'd1;
        12'd414: coeff =  17'd3;
        12'd415: coeff =  17'd1;
        12'd416: coeff = -17'd4;
        12'd417: coeff = -17'd10;
        12'd418: coeff = -17'd11;
        12'd419: coeff = -17'd6;
        12'd420: coeff =  17'd4;
        12'd421: coeff =  17'd15;
        12'd422: coeff =  17'd21;
        12'd423: coeff =  17'd19;
        12'd424: coeff =  17'd8;
        12'd425: coeff = -17'd9;
        12'd426: coeff = -17'd24;
        12'd427: coeff = -17'd31;
        12'd428: coeff = -17'd25;
        12'd429: coeff = -17'd9;
        12'd430: coeff =  17'd13;
        12'd431: coeff =  17'd31;
        12'd432: coeff =  17'd38;
        12'd433: coeff =  17'd29;
        12'd434: coeff =  17'd8;
        12'd435: coeff = -17'd18;
        12'd436: coeff = -17'd37;
        12'd437: coeff = -17'd43;
        12'd438: coeff = -17'd31;
        12'd439: coeff = -17'd6;
        12'd440: coeff =  17'd22;
        12'd441: coeff =  17'd41;
        12'd442: coeff =  17'd44;
        12'd443: coeff =  17'd29;
        12'd444: coeff =  17'd0;
        12'd445: coeff = -17'd30;
        12'd446: coeff = -17'd49;
        12'd447: coeff = -17'd49;
        12'd448: coeff = -17'd29;
        12'd449: coeff =  17'd3;
        12'd450: coeff =  17'd32;
        12'd451: coeff =  17'd45;
        12'd452: coeff =  17'd35;
        12'd453: coeff =  17'd4;
        12'd454: coeff = -17'd37;
        12'd455: coeff = -17'd70;
        12'd456: coeff = -17'd80;
        12'd457: coeff = -17'd61;
        12'd458: coeff = -17'd21;
        12'd459: coeff =  17'd15;
        12'd460: coeff =  17'd20;
        12'd461: coeff = -17'd37;
        12'd462: coeff = -17'd169;
        12'd463: coeff = -17'd373;
        12'd464: coeff =  17'd442;   // This coefficient should be multiplied with the most recent data input
      
        // This should never occur.
        default: coeff =  17'h0000;
      
      endcase
  end

endmodule
